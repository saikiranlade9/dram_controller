`timescale 1 us / 100 ns